----------------------------------------------------------
--	AUTOR: ULISES MARTINEZ RODRIGUEZ
--	DATE: 2020-11-28
--	DESCRIPTION: REALIZA EL DESPLAZAMIENTO DE 1 BIT A
--				LA IZQUIERDA
----------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY BITSHIFT_LEFT_48_BITS IS
	PORT(
		A:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		O:	OUT	STD_LOGIC_VECTOR(47 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE DATAFLOW OF BITSHIFT_LEFT_48_BITS IS
BEGIN
	O(47 DOWNTO 1) <= A(46 DOWNTO 0);
	O(0) <= '0';
END ARCHITECTURE;