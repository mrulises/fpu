----------------------------------------------------------
--	AUTOR: ULISES MARTINEZ RODRIGUEZ
--	DATE: 2020-12-07
--	DESCRIPTION: FUNCION DE EXCEPTION
----------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FUNCTION_E IS
	PORT(
		N, I, S, O, SI:	IN	STD_LOGIC;
		R:				IN	STD_LOGIC_VECTOR(1 DOWNTO 0);
		F:				OUT	STD_LOGIC_VECTOR(31 DOWNTO 0);
		H:				OUT	STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE DATAFLOW OF FUNCTION_E IS

SIGNAL INPUT: STD_LOGIC_VECTOR(6 DOWNTO 0);

BEGIN
	INPUT <= N & I & S & O & R & SI;
	
	F <= SI & "0000000000000000000000000000000" WHEN INPUT(6 DOWNTO 1)="000000" ELSE
		 SI & "1111111111111111111111111111111" WHEN INPUT(6)='1' ELSE
		 SI & "1111111111111111111111111111111" WHEN INPUT(6 DOWNTO 5)="01" ELSE
		 SI & "0000000000000000000000000000000" WHEN INPUT(6 DOWNTO 4)="001" ELSE
		 SI & "1111111011111111111111111111111" WHEN INPUT(6 DOWNTO 1)="000100" ELSE
		 SI & "1111111011111111111111111111111" WHEN INPUT(6 DOWNTO 0)="0001010" ELSE
		 SI & "1111111100000000000000000000000" WHEN INPUT(6 DOWNTO 0)="0001011" ELSE
		 SI & "1111111100000000000000000000000" WHEN INPUT(6 DOWNTO 0)="0001100" ELSE
		 SI & "1111111011111111111111111111111" WHEN INPUT(6 DOWNTO 0)="0001101" ELSE
		 SI & "1111111100000000000000000000000" WHEN INPUT(6 DOWNTO 1)="000111" ELSE
		 SI & "0000000000000000000000000000000";
		 
	H <= "0000" WHEN INPUT(6 DOWNTO 3)="0000" ELSE
		 "1000" WHEN INPUT(6)='1' ELSE
		 "0100" WHEN INPUT(6 DOWNTO 5)="01" ELSE
		 "0010" WHEN INPUT(6 DOWNTO 4)="001" ELSE
		 "0001" WHEN INPUT(6 DOWNTO 3)="0001" ELSE
		 "0000";
		
END ARCHITECTURE;