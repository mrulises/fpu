----------------------------------------------------------
--	AUTOR: ULISES MARTINEZ RODRIGUEZ
--	DATE: 2020-07-12
--	DESCRIPTION: DETERMINA SI ES INFINITO
----------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY IS_INFINITY IS
	PORT(
		I:	IN	STD_LOGIC_VECTOR(30 DOWNTO 0);
		O:	OUT	STD_LOGIC
	);
END ENTITY;

ARCHITECTURE DATAFLOW OF IS_INFINITY IS
BEGIN
	O <= '1' WHEN I="1111111100000000000000000000000" ELSE '0';
END ARCHITECTURE;