----------------------------------------------------------
--	AUTOR: ULISES MARTINEZ RODRIGUEZ
--	DATE: 2020-11-29
--	DESCRIPTION: MULTIPLEXOR DE 128 ENTRADAS A UNA SALIDA
--				DE 96 BITS
----------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MUX_128_TO_1_96_BITS IS
	PORT(
		SEL:	IN	STD_LOGIC_VECTOR(6 DOWNTO 0);
		I_0:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_1:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_2:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_3:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_4:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_5:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_6:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_7:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_8:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_9:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_10:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_11:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_12:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_13:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_14:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_15:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_16:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_17:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_18:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_19:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_20:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_21:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_22:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_23:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_24:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_25:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_26:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_27:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_28:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_29:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_30:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_31:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_32:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_33:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_34:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_35:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_36:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_37:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_38:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_39:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_40:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_41:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_42:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_43:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_44:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_45:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_46:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_47:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_48:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_49:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_50:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_51:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_52:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_53:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_54:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_55:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_56:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_57:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_58:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_59:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_60:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_61:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_62:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_63:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_64:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_65:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_66:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_67:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_68:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_69:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_70:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_71:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_72:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_73:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_74:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_75:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_76:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_77:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_78:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_79:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_80:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_81:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_82:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_83:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_84:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_85:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_86:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_87:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_88:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_89:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_90:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_91:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_92:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_93:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_94:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_95:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_96:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_97:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_98:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_99:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_100:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_101:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_102:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_103:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_104:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_105:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_106:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_107:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_108:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_109:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_110:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_111:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_112:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_113:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_114:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_115:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_116:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_117:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_118:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_119:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_120:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_121:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_122:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_123:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_124:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_125:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_126:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		I_127:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		O:		OUT	STD_LOGIC_VECTOR(95 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE DATAFLOW OF MUX_128_TO_1_96_BITS IS
BEGIN
	WITH SEL SELECT
		O <= I_0 WHEN "0000000",
			I_1 WHEN "0000001",
			I_2 WHEN "0000010",
			I_3 WHEN "0000011",
			I_4 WHEN "0000100",
			I_5 WHEN "0000101",
			I_6 WHEN "0000110",
			I_7 WHEN "0000111",
			I_8 WHEN "0001000",
			I_9 WHEN "0001001",
			I_10 WHEN "0001010",
			I_11 WHEN "0001011",
			I_12 WHEN "0001100",
			I_13 WHEN "0001101",
			I_14 WHEN "0001110",
			I_15 WHEN "0001111",
			I_16 WHEN "0010000",
			I_17 WHEN "0010001",
			I_18 WHEN "0010010",
			I_19 WHEN "0010011",
			I_20 WHEN "0010100",
			I_21 WHEN "0010101",
			I_22 WHEN "0010110",
			I_23 WHEN "0010111",
			I_24 WHEN "0011000",
			I_25 WHEN "0011001",
			I_26 WHEN "0011010",
			I_27 WHEN "0011011",
			I_28 WHEN "0011100",
			I_29 WHEN "0011101",
			I_30 WHEN "0011110",
			I_31 WHEN "0011111",
			I_32 WHEN "0100000",
			I_33 WHEN "0100001",
			I_34 WHEN "0100010",
			I_35 WHEN "0100011",
			I_36 WHEN "0100100",
			I_37 WHEN "0100101",
			I_38 WHEN "0100110",
			I_39 WHEN "0100111",
			I_40 WHEN "0101000",
			I_41 WHEN "0101001",
			I_42 WHEN "0101010",
			I_43 WHEN "0101011",
			I_44 WHEN "0101100",
			I_45 WHEN "0101101",
			I_46 WHEN "0101110",
			I_47 WHEN "0101111",
			I_48 WHEN "0110000",
			I_49 WHEN "0110001",
			I_50 WHEN "0110010",
			I_51 WHEN "0110011",
			I_52 WHEN "0110100",
			I_53 WHEN "0110101",
			I_54 WHEN "0110110",
			I_55 WHEN "0110111",
			I_56 WHEN "0111000",
			I_57 WHEN "0111001",
			I_58 WHEN "0111010",
			I_59 WHEN "0111011",
			I_60 WHEN "0111100",
			I_61 WHEN "0111101",
			I_62 WHEN "0111110",
			I_63 WHEN "0111111",
			I_64 WHEN "1000000",
			I_65 WHEN "1000001",
			I_66 WHEN "1000010",
			I_67 WHEN "1000011",
			I_68 WHEN "1000100",
			I_69 WHEN "1000101",
			I_70 WHEN "1000110",
			I_71 WHEN "1000111",
			I_72 WHEN "1001000",
			I_73 WHEN "1001001",
			I_74 WHEN "1001010",
			I_75 WHEN "1001011",
			I_76 WHEN "1001100",
			I_77 WHEN "1001101",
			I_78 WHEN "1001110",
			I_79 WHEN "1001111",
			I_80 WHEN "1010000",
			I_81 WHEN "1010001",
			I_82 WHEN "1010010",
			I_83 WHEN "1010011",
			I_84 WHEN "1010100",
			I_85 WHEN "1010101",
			I_86 WHEN "1010110",
			I_87 WHEN "1010111",
			I_88 WHEN "1011000",
			I_89 WHEN "1011001",
			I_90 WHEN "1011010",
			I_91 WHEN "1011011",
			I_92 WHEN "1011100",
			I_93 WHEN "1011101",
			I_94 WHEN "1011110",
			I_95 WHEN "1011111",
			I_96 WHEN "1100000",
			I_97 WHEN "1100001",
			I_98 WHEN "1100010",
			I_99 WHEN "1100011",
			I_100 WHEN "1100100",
			I_101 WHEN "1100101",
			I_102 WHEN "1100110",
			I_103 WHEN "1100111",
			I_104 WHEN "1101000",
			I_105 WHEN "1101001",
			I_106 WHEN "1101010",
			I_107 WHEN "1101011",
			I_108 WHEN "1101100",
			I_109 WHEN "1101101",
			I_110 WHEN "1101110",
			I_111 WHEN "1101111",
			I_112 WHEN "1110000",
			I_113 WHEN "1110001",
			I_114 WHEN "1110010",
			I_115 WHEN "1110011",
			I_116 WHEN "1110100",
			I_117 WHEN "1110101",
			I_118 WHEN "1110110",
			I_119 WHEN "1110111",
			I_120 WHEN "1111000",
			I_121 WHEN "1111001",
			I_122 WHEN "1111010",
			I_123 WHEN "1111011",
			I_124 WHEN "1111100",
			I_125 WHEN "1111101",
			I_126 WHEN "1111110",
			I_127 WHEN OTHERS;
END ARCHITECTURE;