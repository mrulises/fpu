----------------------------------------------------------
--	AUTOR: ULISES MARTINEZ RODRIGUEZ
--	DATE: 2020-11-29
--	DESCRIPTION: UNIDAD DE PUNTO FLOTANTE PARA PRODUCTO
----------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FPU IS
	PORT(
		A:	IN	STD_LOGIC_VECTOR(31 DOWNTO 0);
		B:	IN	STD_LOGIC_VECTOR(31 DOWNTO 0);
		R:	IN	STD_LOGIC_VECTOR(1 DOWNTO 0);
		C:	OUT	STD_LOGIC_VECTOR(31 DOWNTO 0);
		H:	OUT	STD_LOGIC_VECTOR(2 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE STRUCUTURE OF FPU IS

COMPONENT XOR_C IS
	PORT(
		X:		IN		STD_LOGIC;
		Y:		IN		STD_LOGIC;
		Z:		OUT		STD_LOGIC
	);
END COMPONENT;

COMPONENT ADD_10_BITS IS
	PORT(
		CARRYIN:	IN	STD_LOGIC;
		ADDEND1:	IN	STD_LOGIC_VECTOR(9 DOWNTO 0);
		ADDEND2:	IN	STD_LOGIC_VECTOR(9 DOWNTO 0);
		SUM:		OUT	STD_LOGIC_VECTOR(9 DOWNTO 0);
		CARRYOUT:	OUT	STD_LOGIC
	);
END COMPONENT;

COMPONENT MUX_2_TO_1_10_BITS IS
	PORT(
		SEL:	IN	STD_LOGIC;
		I_0:	IN	STD_LOGIC_VECTOR(9 DOWNTO 0);
		I_1:	IN	STD_LOGIC_VECTOR(9 DOWNTO 0);
		O:		OUT	STD_LOGIC_VECTOR(9 DOWNTO 0)
	);
END COMPONENT;

COMPONENT RECOVER_BIT IS
	PORT(
		E:		IN	STD_LOGIC_VECTOR(7 DOWNTO 0);
		M:		IN 	STD_LOGIC_VECTOR(22 DOWNTO 0);
		P:		OUT	STD_LOGIC_VECTOR(23 DOWNTO 0)
	);
END COMPONENT;

COMPONENT MULT_24_BITS IS
	PORT(
		MULTIPLICAND:	IN	STD_LOGIC_VECTOR(23 DOWNTO 0);
		MULTIPLIER:		IN	STD_LOGIC_VECTOR(23 DOWNTO 0);
		PRODUCTHIGH:	OUT	STD_LOGIC_VECTOR(23 DOWNTO 0);
		PRODUCTLOW:		OUT	STD_LOGIC_VECTOR(23 DOWNTO 0)
	);
END COMPONENT;

COMPONENT FORMAT_MULT IS
	PORT(
		H:		IN	STD_LOGIC_VECTOR(23 DOWNTO 0);
		L:		IN	STD_LOGIC_VECTOR(23 DOWNTO 0);
		M:		OUT	STD_LOGIC_VECTOR(47 DOWNTO 0)
	);
END COMPONENT;

COMPONENT NORMALIZER IS
	PORT(
		S:		IN	STD_LOGIC;
		E:		IN	STD_LOGIC_VECTOR(9 DOWNTO 0);
		M:		IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		OS:		OUT	STD_LOGIC;
		OE:		OUT	STD_LOGIC_VECTOR(9 DOWNTO 0);
		OM:		OUT	STD_LOGIC_VECTOR(47 DOWNTO 0)
	);
END COMPONENT;

COMPONENT ROUND IS
	PORT(
		R:	IN	STD_LOGIC_VECTOR(1 DOWNTO 0);
		S:	IN	STD_LOGIC;
		E:	IN	STD_LOGIC_VECTOR(9 DOWNTO 0);
		M:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		F:	OUT	STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

SIGNAL NORMA_S:		STD_LOGIC;
SIGNAL NORMA_E:		STD_LOGIC_VECTOR(9 DOWNTO 0);
SIGNAL REGISTER_B:	STD_LOGIC_VECTOR(9 DOWNTO 0):="0100000001";
SIGNAL REGISTER_O:	STD_LOGIC_VECTOR(9 DOWNTO 0):="0000000001";
SIGNAL ADD_INP_A:	STD_LOGIC_VECTOR(9 DOWNTO 0);
SIGNAL ADD_MUX_A:	STD_LOGIC_VECTOR(9 DOWNTO 0);
SIGNAL ADD_MUX_B:	STD_LOGIC_VECTOR(9 DOWNTO 0);
SIGNAL MULT_INP_A:	STD_LOGIC_VECTOR(23 DOWNTO 0);
SIGNAL MULT_INP_B:	STD_LOGIC_VECTOR(23 DOWNTO 0);
SIGNAL MULT_R_H:	STD_LOGIC_VECTOR(23 DOWNTO 0);
SIGNAL MULT_R_L:	STD_LOGIC_VECTOR(23 DOWNTO 0);
SIGNAL NORMA_M:		STD_LOGIC_VECTOR(47 DOWNTO 0);
SIGNAL O_NORMA_S:	STD_LOGIC;
SIGNAL O_NORMA_E:	STD_LOGIC_VECTOR(9 DOWNTO 0);
SIGNAL O_NORMA_M:	STD_LOGIC_VECTOR(47 DOWNTO 0);
SIGNAL F:			STD_LOGIC_VECTOR(31 DOWNTO 0);

BEGIN
	
	C_XOR_C:	XOR_C PORT MAP(A(31), B(31), NORMA_S);
	ADD_B:		ADD_10_BITS PORT MAP('0', ADD_MUX_A, REGISTER_B, ADD_INP_A, OPEN);
	ADD_E:		ADD_10_BITS PORT MAP('0', ADD_INP_A, ADD_MUX_B, NORMA_E, OPEN);
	RECOVER_A:	RECOVER_BIT PORT MAP(A(30 DOWNTO 23), A(22 DOWNTO 0), MULT_INP_A);
	RECOVER_B:	RECOVER_BIT PORT MAP(B(30 DOWNTO 23), B(22 DOWNTO 0), MULT_INP_B);
	MULT:		MULT_24_BITS PORT MAP(MULT_INP_A, MULT_INP_B, MULT_R_H, MULT_R_L);
	FORMAT:		FORMAT_MULT PORT MAP(MULT_R_H, MULT_R_L, NORMA_M);
	NORMA:		NORMALIZER PORT MAP(NORMA_S, NORMA_E, NORMA_M, O_NORMA_S, O_NORMA_E, O_NORMA_M);
	MUX_A:		MUX_2_TO_1_10_BITS PORT MAP(MULT_INP_A(23), REGISTER_O, "00" & A(30 DOWNTO 23), ADD_MUX_A);
	MUX_B:		MUX_2_TO_1_10_BITS PORT MAP(MULT_INP_B(23), REGISTER_O, "00" & B(30 DOWNTO 23), ADD_MUX_B);
	ROUN:		ROUND PORT MAP(R, O_NORMA_S, O_NORMA_E, O_NORMA_M, F);
	
	C <= F;
	
END ARCHITECTURE;