----------------------------------------------------------
--	AUTOR: ULISES MARTINEZ RODRIGUEZ
--	DATE: 2020-11-28
--	DESCRIPTION: MULTIPLEXOR DE 2 ENTRADAS A UNA SALIDA
--				DE 1O BITS
----------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MUX_2_TO_1_10_BITS IS
	PORT(
		SEL:	IN	STD_LOGIC;
		I_0:	IN	STD_LOGIC_VECTOR(9 DOWNTO 0);
		I_1:	IN	STD_LOGIC_VECTOR(9 DOWNTO 0);
		O:		OUT	STD_LOGIC_VECTOR(9 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE DATAFLOW OF MUX_2_TO_1_10_BITS IS
BEGIN
	WITH SEL SELECT
		O	<=	I_0 WHEN '0',
				I_1 WHEN OTHERS;
END ARCHITECTURE;