----------------------------------------------------------
--	AUTOR: ULISES MARTINEZ RODRIGUEZ
--	DATE: 2020-11-28
--	DESCRIPTION: MULTIPLEXOR DE 64 ENTRADAS A UNA SALIDA
--				DE 48 BITS
----------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MUX_64_TO_1_48_BITS IS
	PORT(
		SEL:	IN	STD_LOGIC_VECTOR(5 DOWNTO 0);
		I_0:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_1:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_2:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_3:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_4:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_5:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_6:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_7:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_8:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_9:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_10:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_11:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_12:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_13:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_14:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_15:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_16:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_17:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_18:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_19:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_20:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_21:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_22:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_23:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_24:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_25:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_26:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_27:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_28:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_29:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_30:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_31:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_32:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_33:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_34:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_35:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_36:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_37:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_38:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_39:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_40:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_41:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_42:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_43:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_44:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_45:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_46:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_47:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_48:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_49:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_50:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_51:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_52:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_53:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_54:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_55:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_56:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_57:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_58:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_59:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_60:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_61:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_62:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_63:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		O:		OUT	STD_LOGIC_VECTOR(47 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE DATAFLOW OF MUX_64_TO_1_48_BITS IS
BEGIN
	WITH SEL SELECT
		O	<=	I_0 WHEN "000000",
			I_1 WHEN "000001",
			I_2 WHEN "000010",
			I_3 WHEN "000011",
			I_4 WHEN "000100",
			I_5 WHEN "000101",
			I_6 WHEN "000110",
			I_7 WHEN "000111",
			I_8 WHEN "001000",
			I_9 WHEN "001001",
			I_10 WHEN "001010",
			I_11 WHEN "001011",
			I_12 WHEN "001100",
			I_13 WHEN "001101",
			I_14 WHEN "001110",
			I_15 WHEN "001111",
			I_16 WHEN "010000",
			I_17 WHEN "010001",
			I_18 WHEN "010010",
			I_19 WHEN "010011",
			I_20 WHEN "010100",
			I_21 WHEN "010101",
			I_22 WHEN "010110",
			I_23 WHEN "010111",
			I_24 WHEN "011000",
			I_25 WHEN "011001",
			I_26 WHEN "011010",
			I_27 WHEN "011011",
			I_28 WHEN "011100",
			I_29 WHEN "011101",
			I_30 WHEN "011110",
			I_31 WHEN "011111",
			I_32 WHEN "100000",
			I_33 WHEN "100001",
			I_34 WHEN "100010",
			I_35 WHEN "100011",
			I_36 WHEN "100100",
			I_37 WHEN "100101",
			I_38 WHEN "100110",
			I_39 WHEN "100111",
			I_40 WHEN "101000",
			I_41 WHEN "101001",
			I_42 WHEN "101010",
			I_43 WHEN "101011",
			I_44 WHEN "101100",
			I_45 WHEN "101101",
			I_46 WHEN "101110",
			I_47 WHEN "101111",
			I_48 WHEN "110000",
			I_49 WHEN "110001",
			I_50 WHEN "110010",
			I_51 WHEN "110011",
			I_52 WHEN "110100",
			I_53 WHEN "110101",
			I_54 WHEN "110110",
			I_55 WHEN "110111",
			I_56 WHEN "111000",
			I_57 WHEN "111001",
			I_58 WHEN "111010",
			I_59 WHEN "111011",
			I_60 WHEN "111100",
			I_61 WHEN "111101",
			I_62 WHEN "111110",
			I_63 WHEN OTHERS;
END ARCHITECTURE;