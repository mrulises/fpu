----------------------------------------------------------
--	AUTOR: ULISES MARTINEZ RODRIGUEZ
--	DATE: 2020-11-28
--	DESCRIPTION: REALIZA UN COMPLEMENTO A DOS DEL LA
--				ENTRADA
----------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY TWO_S_COMPLE_10_BITS IS
	PORT(
		A:		IN	STD_LOGIC_VECTOR(9 DOWNTO 0);
		C:		OUT	STD_LOGIC_VECTOR(9 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE STRUCTURE OF TWO_S_COMPLE_10_BITS IS

COMPONENT ADD_10_BITS IS
	PORT(
		CARRYIN:	IN	STD_LOGIC;
		ADDEND1:	IN	STD_LOGIC_VECTOR(9 DOWNTO 0);
		ADDEND2:	IN	STD_LOGIC_VECTOR(9 DOWNTO 0);
		SUM:		OUT	STD_LOGIC_VECTOR(9 DOWNTO 0);
		CARRYOUT:	OUT	STD_LOGIC
	);
END COMPONENT;

COMPONENT NOT_10_BITS IS
	PORT(
		I:	IN	STD_LOGIC_VECTOR(9 DOWNTO 0);
		O:	OUT	STD_LOGIC_VECTOR(9 DOWNTO 0)
	);
END COMPONENT;

SIGNAL COMPLEMENT:		STD_LOGIC_VECTOR(9 DOWNTO 0);

BEGIN
	
	NOT_C:	NOT_10_BITS PORT MAP(A, COMPLEMENT);
	COMPLEMENT2:	ADD_10_BITS PORT MAP('0', COMPLEMENT, "0000000001", C, OPEN);
	
END ARCHITECTURE;