----------------------------------------------------------
--	AUTOR: ULISES MARTINEZ RODRIGUEZ
--	DATE: 2020-11-28
--	DESCRIPTION: NORMALIZA UN NUMERO DE PUNTO FLOTANTE
----------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY NORMALIZER IS
	PORT(
		S:		IN	STD_LOGIC;
		E:		IN	STD_LOGIC_VECTOR(9 DOWNTO 0);
		M:		IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		OS:		OUT	STD_LOGIC;
		OE:		OUT	STD_LOGIC_VECTOR(9 DOWNTO 0);
		OM:		OUT	STD_LOGIC_VECTOR(47 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE STRUCTURE OF NORMALIZER IS

COMPONENT FUNCTION_D IS
	PORT(
		M:		IN	STD_LOGIC_VECTOR(46 DOWNTO 0);
		POSS:	OUT	STD_LOGIC_VECTOR(5 DOWNTO 0)
	);
END COMPONENT;

COMPONENT TWO_S_COMPLE_10_BITS IS
	PORT(
		A:		IN	STD_LOGIC_VECTOR(9 DOWNTO 0);
		C:		OUT	STD_LOGIC_VECTOR(9 DOWNTO 0)
	);
END COMPONENT;

COMPONENT ADD_10_BITS IS
	PORT(
		CARRYIN:	IN	STD_LOGIC;
		ADDEND1:	IN	STD_LOGIC_VECTOR(9 DOWNTO 0);
		ADDEND2:	IN	STD_LOGIC_VECTOR(9 DOWNTO 0);
		SUM:		OUT	STD_LOGIC_VECTOR(9 DOWNTO 0);
		CARRYOUT:	OUT	STD_LOGIC
	);
END COMPONENT;

COMPONENT MUX_2_TO_1_10_BITS IS
	PORT(
		SEL:	IN	STD_LOGIC;
		I_0:	IN	STD_LOGIC_VECTOR(9 DOWNTO 0);
		I_1:	IN	STD_LOGIC_VECTOR(9 DOWNTO 0);
		O:		OUT	STD_LOGIC_VECTOR(9 DOWNTO 0)
	);
END COMPONENT;

COMPONENT MUX_2_TO_1_48_BITS IS
	PORT(
		SEL:	IN	STD_LOGIC;
		I_0:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_1:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		O:		OUT	STD_LOGIC_VECTOR(47 DOWNTO 0)
	);
END COMPONENT;

COMPONENT MUX_64_TO_1_48_BITS IS
	PORT(
		SEL:	IN	STD_LOGIC_VECTOR(5 DOWNTO 0);
		I_0:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_1:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_2:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_3:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_4:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_5:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_6:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_7:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_8:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_9:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_10:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_11:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_12:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_13:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_14:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_15:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_16:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_17:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_18:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_19:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_20:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_21:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_22:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_23:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_24:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_25:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_26:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_27:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_28:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_29:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_30:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_31:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_32:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_33:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_34:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_35:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_36:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_37:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_38:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_39:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_40:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_41:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_42:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_43:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_44:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_45:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_46:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_47:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_48:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_49:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_50:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_51:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_52:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_53:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_54:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_55:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_56:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_57:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_58:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_59:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_60:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_61:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_62:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		I_63:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		O:		OUT	STD_LOGIC_VECTOR(47 DOWNTO 0)
	);
END COMPONENT;

COMPONENT BITSHIFT_LEFT_48_BITS IS
	PORT(
		A:	IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
		O:	OUT	STD_LOGIC_VECTOR(47 DOWNTO 0)
	);
END COMPONENT;

SIGNAL O_FUNCTION_D:	STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL O_TWO_S:			STD_LOGIC_VECTOR(9 DOWNTO 0);
SIGNAL REGISTER_1:		STD_LOGIC_VECTOR(9 DOWNTO 0):= "0000000001";
SIGNAL O_MUX_E:			STD_LOGIC_VECTOR(9 DOWNTO 0);
SIGNAL O_MUX_S:			STD_LOGIC_VECTOR(47 DOWNTO 0);
SIGNAL BS_R:			STD_LOGIC_VECTOR(2255 DOWNTO 0);

BEGIN
	
	E_FUNCTION_D:	FUNCTION_D PORT MAP(M(46 DOWNTO 0), O_FUNCTION_D);
	E_TWO_S:		TWO_S_COMPLE_10_BITS PORT MAP("0000" & O_FUNCTION_D, O_TWO_S);
	MUX_E:			MUX_2_TO_1_10_BITS PORT MAP(M(47), O_TWO_S, REGISTER_1, O_MUX_E);
	ADD:			ADD_10_BITS PORT MAP('0', E, O_MUX_E, OE, OPEN);
	MUX_M:			MUX_2_TO_1_48_BITS PORT MAP(M(47), O_MUX_S, M, OM);
	BS1:			BITSHIFT_LEFT_48_BITS PORT MAP(M, BS_R(47 DOWNTO 0));
	BS2:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(47 DOWNTO 0), BS_R(95 DOWNTO 48));
	BS3:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(95 DOWNTO 48), BS_R(143 DOWNTO 96));
	BS4:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(143 DOWNTO 96), BS_R(191 DOWNTO 144));
	BS5:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(191 DOWNTO 144), BS_R(239 DOWNTO 192));
	BS6:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(239 DOWNTO 192), BS_R(287 DOWNTO 240));
	BS7:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(287 DOWNTO 240), BS_R(335 DOWNTO 288));
	BS8:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(335 DOWNTO 288), BS_R(383 DOWNTO 336));
	BS9:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(383 DOWNTO 336), BS_R(431 DOWNTO 384));
	BS10:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(431 DOWNTO 384), BS_R(479 DOWNTO 432));
	BS11:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(479 DOWNTO 432), BS_R(527 DOWNTO 480));
	BS12:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(527 DOWNTO 480), BS_R(575 DOWNTO 528));
	BS13:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(575 DOWNTO 528), BS_R(623 DOWNTO 576));
	BS14:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(623 DOWNTO 576), BS_R(671 DOWNTO 624));
	BS15:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(671 DOWNTO 624), BS_R(719 DOWNTO 672));
	BS16:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(719 DOWNTO 672), BS_R(767 DOWNTO 720));
	BS17:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(767 DOWNTO 720), BS_R(815 DOWNTO 768));
	BS18:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(815 DOWNTO 768), BS_R(863 DOWNTO 816));
	BS19:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(863 DOWNTO 816), BS_R(911 DOWNTO 864));
	BS20:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(911 DOWNTO 864), BS_R(959 DOWNTO 912));
	BS21:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(959 DOWNTO 912), BS_R(1007 DOWNTO 960));
	BS22:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(1007 DOWNTO 960), BS_R(1055 DOWNTO 1008));
	BS23:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(1055 DOWNTO 1008), BS_R(1103 DOWNTO 1056));
	BS24:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(1103 DOWNTO 1056), BS_R(1151 DOWNTO 1104));
	BS25:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(1151 DOWNTO 1104), BS_R(1199 DOWNTO 1152));
	BS26:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(1199 DOWNTO 1152), BS_R(1247 DOWNTO 1200));
	BS27:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(1247 DOWNTO 1200), BS_R(1295 DOWNTO 1248));
	BS28:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(1295 DOWNTO 1248), BS_R(1343 DOWNTO 1296));
	BS29:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(1343 DOWNTO 1296), BS_R(1391 DOWNTO 1344));
	BS30:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(1391 DOWNTO 1344), BS_R(1439 DOWNTO 1392));
	BS31:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(1439 DOWNTO 1392), BS_R(1487 DOWNTO 1440));
	BS32:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(1487 DOWNTO 1440), BS_R(1535 DOWNTO 1488));
	BS33:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(1535 DOWNTO 1488), BS_R(1583 DOWNTO 1536));
	BS34:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(1583 DOWNTO 1536), BS_R(1631 DOWNTO 1584));
	BS35:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(1631 DOWNTO 1584), BS_R(1679 DOWNTO 1632));
	BS36:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(1679 DOWNTO 1632), BS_R(1727 DOWNTO 1680));
	BS37:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(1727 DOWNTO 1680), BS_R(1775 DOWNTO 1728));
	BS38:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(1775 DOWNTO 1728), BS_R(1823 DOWNTO 1776));
	BS39:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(1823 DOWNTO 1776), BS_R(1871 DOWNTO 1824));
	BS40:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(1871 DOWNTO 1824), BS_R(1919 DOWNTO 1872));
	BS41:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(1919 DOWNTO 1872), BS_R(1967 DOWNTO 1920));
	BS42:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(1967 DOWNTO 1920), BS_R(2015 DOWNTO 1968));
	BS43:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(2015 DOWNTO 1968), BS_R(2063 DOWNTO 2016));
	BS44:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(2063 DOWNTO 2016), BS_R(2111 DOWNTO 2064));
	BS45:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(2111 DOWNTO 2064), BS_R(2159 DOWNTO 2112));
	BS46:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(2159 DOWNTO 2112), BS_R(2207 DOWNTO 2160));
	BS47:			BITSHIFT_LEFT_48_BITS PORT MAP(BS_R(2207 DOWNTO 2160), BS_R(2255 DOWNTO 2208));
	MUX_S:			MUX_64_TO_1_48_BITS PORT MAP(O_FUNCTION_D, BS_R(47 DOWNTO 0), BS_R(95 DOWNTO 48), BS_R(143 DOWNTO 96), BS_R(191 DOWNTO 144), BS_R(239 DOWNTO 192), BS_R(287 DOWNTO 240), BS_R(335 DOWNTO 288), BS_R(383 DOWNTO 336), BS_R(431 DOWNTO 384), BS_R(479 DOWNTO 432), BS_R(527 DOWNTO 480), 
					BS_R(575 DOWNTO 528), BS_R(623 DOWNTO 576), BS_R(671 DOWNTO 624), BS_R(719 DOWNTO 672), BS_R(767 DOWNTO 720), BS_R(815 DOWNTO 768), BS_R(863 DOWNTO 816), BS_R(911 DOWNTO 864), BS_R(959 DOWNTO 912), BS_R(1007 DOWNTO 960), 
					BS_R(1055 DOWNTO 1008), BS_R(1103 DOWNTO 1056), BS_R(1151 DOWNTO 1104), BS_R(1199 DOWNTO 1152), BS_R(1247 DOWNTO 1200), BS_R(1295 DOWNTO 1248), BS_R(1343 DOWNTO 1296), BS_R(1391 DOWNTO 1344), BS_R(1439 DOWNTO 1392), BS_R(1487 DOWNTO 1440), 
					BS_R(1535 DOWNTO 1488), BS_R(1583 DOWNTO 1536), BS_R(1631 DOWNTO 1584), BS_R(1679 DOWNTO 1632), BS_R(1727 DOWNTO 1680), BS_R(1775 DOWNTO 1728), BS_R(1823 DOWNTO 1776), BS_R(1871 DOWNTO 1824), BS_R(1919 DOWNTO 1872), BS_R(1967 DOWNTO 1920), 
					BS_R(2015 DOWNTO 1968), BS_R(2063 DOWNTO 2016), BS_R(2111 DOWNTO 2064), BS_R(2159 DOWNTO 2112), BS_R(2207 DOWNTO 2160), BS_R(2255 DOWNTO 2208), "000000000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000000000", 
					"000000000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000000000", 
					"000000000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000000000", "000000000000000000000000000000000000000000000000", O_MUX_S);
	OS <= S;
	
END ARCHITECTURE;