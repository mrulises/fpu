----------------------------------------------------------
--	AUTOR: ULISES MARTINEZ RODRIGUEZ
--	DATE: 2020-11-28
--	DESCRIPTION: FUNCION PARA DETERMINAR LA POSICION DEL
--				BIT MAS SIGNIFICATIVO EN 1
----------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FUNCTION_D IS
	PORT(
		M:		IN	STD_LOGIC_VECTOR(46 DOWNTO 0);
		POSS:	OUT	STD_LOGIC_VECTOR(5 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE DATAFLOW OF FUNCTION_D IS
BEGIN
	POSS <= "000000" WHEN M(46)='1' ELSE
			"000001" WHEN M(45)='1' ELSE
			"000010" WHEN M(44)='1' ELSE
			"000011" WHEN M(43)='1' ELSE
			"000100" WHEN M(42)='1' ELSE
			"000101" WHEN M(41)='1' ELSE
			"000110" WHEN M(40)='1' ELSE
			"000111" WHEN M(39)='1' ELSE
			"001000" WHEN M(38)='1' ELSE
			"001001" WHEN M(37)='1' ELSE
			"001010" WHEN M(36)='1' ELSE
			"001011" WHEN M(35)='1' ELSE
			"001100" WHEN M(34)='1' ELSE
			"001101" WHEN M(33)='1' ELSE
			"001110" WHEN M(32)='1' ELSE
			"001111" WHEN M(31)='1' ELSE
			"010000" WHEN M(30)='1' ELSE
			"010001" WHEN M(29)='1' ELSE
			"010010" WHEN M(28)='1' ELSE
			"010011" WHEN M(27)='1' ELSE
			"010100" WHEN M(26)='1' ELSE
			"010101" WHEN M(25)='1' ELSE
			"010110" WHEN M(24)='1' ELSE
			"010111" WHEN M(23)='1' ELSE
			"011000" WHEN M(22)='1' ELSE
			"011001" WHEN M(21)='1' ELSE
			"011010" WHEN M(20)='1' ELSE
			"011011" WHEN M(19)='1' ELSE
			"011100" WHEN M(18)='1' ELSE
			"011101" WHEN M(17)='1' ELSE
			"011110" WHEN M(16)='1' ELSE
			"011111" WHEN M(15)='1' ELSE
			"100000" WHEN M(14)='1' ELSE
			"100001" WHEN M(13)='1' ELSE
			"100010" WHEN M(12)='1' ELSE
			"100011" WHEN M(11)='1' ELSE
			"100100" WHEN M(10)='1' ELSE
			"100101" WHEN M(9)='1' ELSE
			"100110" WHEN M(8)='1' ELSE
			"100111" WHEN M(7)='1' ELSE
			"101000" WHEN M(6)='1' ELSE
			"101001" WHEN M(5)='1' ELSE
			"101010" WHEN M(4)='1' ELSE
			"101011" WHEN M(3)='1' ELSE
			"101100" WHEN M(2)='1' ELSE
			"101101" WHEN M(1)='1' ELSE
			"101110" WHEN M(0)='1' ELSE
			"111111";

END ARCHITECTURE;