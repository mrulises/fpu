----------------------------------------------------------
--	AUTOR: ULISES MARTINEZ RODRIGUEZ
--	DATE: 2020-11-26
--	DESCRIPTION: FORMATEA EL RESULTADO DE UN PRODUCTO
--				DE 24 BITS
----------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FORMAT_MULT IS
	PORT(
		H:		IN	STD_LOGIC_VECTOR(23 DOWNTO 0);
		L:		IN	STD_LOGIC_VECTOR(23 DOWNTO 0);
		M:		OUT	STD_LOGIC_VECTOR(47 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE DATAFLOW OF FORMAT_MULT IS
BEGIN
	M(47 DOWNTO 24) <= H;
	M(23 DOWNTO 0) <= L;
END ARCHITECTURE;