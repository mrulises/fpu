------------------------------------------------
--	AUTOR: ULISES MARTINEZ RODRIGUEZ
--	DATE: 2020-11-25
--	DESCRIPTION: SUMA DE DOS ENTRADAS DE 10 BITS
------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ADD_10_BITS IS
	PORT(
		CARRYIN:	IN	STD_LOGIC;
		ADDEND1:	IN	STD_LOGIC_VECTOR(9 DOWNTO 0);
		ADDEND2:	IN	STD_LOGIC_VECTOR(9 DOWNTO 0);
		SUM:		OUT	STD_LOGIC_VECTOR(9 DOWNTO 0);
		CARRYOUT:	OUT	STD_LOGIC
	);
END ENTITY;

ARCHITECTURE DATAFLOW OF ADD_10_BITS IS

SIGNAL	CARRIES:		STD_LOGIC_VECTOR(10 DOWNTO 0);

	BEGIN
		CARRIES(0) <= CARRYIN;
		
		SUM(0) <= (ADDEND1(0) XOR ADDEND2(0)) XOR CARRIES(0);
		CARRIES(1) <= (ADDEND1(0) AND ADDEND2(0)) OR ((ADDEND1(0) OR ADDEND2(0)) AND CARRIES(0));
		
		SUM(1) <= (ADDEND1(1) XOR ADDEND2(1)) XOR CARRIES(1);
		CARRIES(2) <= (ADDEND1(1) AND ADDEND2(1)) OR ((ADDEND1(1) OR ADDEND2(1)) AND CARRIES(1));
		
		SUM(2) <= (ADDEND1(2) XOR ADDEND2(2)) XOR CARRIES(2);
		CARRIES(3) <= (ADDEND1(2) AND ADDEND2(2)) OR ((ADDEND1(2) OR ADDEND2(2)) AND CARRIES(2));
		
		SUM(3) <= (ADDEND1(3) XOR ADDEND2(3)) XOR CARRIES(3);
		CARRIES(4) <= (ADDEND1(3) AND ADDEND2(3)) OR ((ADDEND1(3) OR ADDEND2(3)) AND CARRIES(3));
		
		SUM(4) <= (ADDEND1(4) XOR ADDEND2(4)) XOR CARRIES(4);
		CARRIES(5) <= (ADDEND1(4) AND ADDEND2(4)) OR ((ADDEND1(4) OR ADDEND2(4)) AND CARRIES(4));
		
		SUM(5) <= (ADDEND1(5) XOR ADDEND2(5)) XOR CARRIES(5);		
		CARRIES(6) <= (ADDEND1(5) AND ADDEND2(5)) OR ((ADDEND1(5) OR ADDEND2(5)) AND CARRIES(5));
		
		SUM(6) <= (ADDEND1(6) XOR ADDEND2(6)) XOR CARRIES(6);
		CARRIES(7) <= (ADDEND1(6) AND ADDEND2(6)) OR ((ADDEND1(6) OR ADDEND2(6)) AND CARRIES(6));
		
		SUM(7) <= (ADDEND1(7) XOR ADDEND2(7)) XOR CARRIES(7);
		CARRIES(8) <= (ADDEND1(7) AND ADDEND2(7)) OR ((ADDEND1(7) OR ADDEND2(7)) AND CARRIES(7));
		
		SUM(8) <= (ADDEND1(8) XOR ADDEND2(8)) XOR CARRIES(8);
		CARRIES(9) <= (ADDEND1(8) AND ADDEND2(8)) OR ((ADDEND1(8) OR ADDEND2(8)) AND CARRIES(8));
		
		SUM(9) <= (ADDEND1(9) XOR ADDEND2(9)) XOR CARRIES(9);
		CARRIES(10) <= (ADDEND1(9) AND ADDEND2(9)) OR ((ADDEND1(9) OR ADDEND2(9)) AND CARRIES(9));
		
		CARRYOUT <= CARRIES(10);
END ARCHITECTURE;