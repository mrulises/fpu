----------------------------------------------------------
--	AUTOR: ULISES MARTINEZ RODRIGUEZ
--	DATE: 2020-11-29
--	DESCRIPTION: DETERMINAR SI SE SUMA 1 PARA EL REDONDEO
----------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FUNCTION_R IS
	PORT(
		R:	IN	STD_LOGIC_VECTOR(1 DOWNTO 0);
		S:	IN	STD_LOGIC;
		RT:	IN	STD_LOGIC;
		ST:	IN	STD_LOGIC;
		V:	OUT	STD_LOGIC
	);
END ENTITY;

ARCHITECTURE DATAFLOW OF FUNCTION_R IS

SIGNAL REG:	STD_LOGIC_VECTOR(4 DOWNTO 0);

BEGIN
	
	REG(4 DOWNTO 3) <= R;
	REG(2) <= S;
	REG(1) <= RT;
	REG(0) <= ST;
	
	V	<= 	'0' WHEN REG(4 DOWNTO 3)="00" ELSE
			'0' WHEN REG(4 DOWNTO 2)="010" ELSE
			'0' WHEN REG(4 DOWNTO 0)="01100" ELSE
			'1' WHEN REG(4 DOWNTO 0)="01101" ELSE
			'1' WHEN REG(4 DOWNTO 0)="01110" ELSE
			'1' WHEN REG(4 DOWNTO 0)="01111" ELSE
			'0' WHEN REG(4 DOWNTO 0)="10000" ELSE
			'1' WHEN REG(4 DOWNTO 0)="10001" ELSE
			'1' WHEN REG(4 DOWNTO 0)="10010" ELSE
			'1' WHEN REG(4 DOWNTO 0)="10011" ELSE
			'0' WHEN REG(4 DOWNTO 2)="101" ELSE
			'0' WHEN REG(4 DOWNTO 0)="11000" ELSE
			'0' WHEN REG(4 DOWNTO 0)="11001" ELSE
			'0' WHEN REG(4 DOWNTO 0)="11010" ELSE
			'1' WHEN REG(4 DOWNTO 0)="11011" ELSE
			'0' WHEN REG(4 DOWNTO 0)="11100" ELSE
			'0' WHEN REG(4 DOWNTO 0)="11101" ELSE
			'0' WHEN REG(4 DOWNTO 0)="11110" ELSE
			'1' WHEN REG(4 DOWNTO 0)="11111" ELSE
			'0';
	
END ARCHITECTURE;