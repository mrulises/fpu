----------------------------------------------------------
--	AUTOR: ULISES MARTINEZ RODRIGUEZ
--	DATE: 2020-07-12
--	DESCRIPTION: DETERMINA SI ES ZERO
----------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY IS_ZERO IS
	PORT(
		I:	IN	STD_LOGIC_VECTOR(30 DOWNTO 0);
		O:	OUT	STD_LOGIC
	);
END ENTITY;

ARCHITECTURE DATAFLOW OF IS_ZERO IS
BEGIN
	O <= NOT( I(30) OR I(29) OR I(28) OR I(27) OR I(26) OR I(25) OR I(24) OR I(23) OR I(22) OR I(21) OR I(20) OR I(19) OR I(18) OR I(17) OR I(16) OR I(15) OR I(14) OR I(13) OR I(12) OR I(11) OR I(10) OR I(9) OR I(8) OR I(7) OR I(6) OR I(5) OR I(4) OR I(3) OR I(2) OR I(1) OR I(0));
END ARCHITECTURE;