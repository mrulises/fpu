----------------------------------------------------------
--	AUTOR: ULISES MARTINEZ RODRIGUEZ
--	DATE: 2020-12-07
--	DESCRIPTION: GENERADOR DE EXCEPCIONES
----------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY EXCEPTIONS IS
	PORT(
		A:		IN	STD_LOGIC_VECTOR(31 DOWNTO 0);
		B:		IN	STD_LOGIC_VECTOR(31 DOWNTO 0);
		C:		IN	STD_LOGIC_VECTOR(31 DOWNTO 0);
		R:		IN	STD_LOGIC_VECTOR(1 DOWNTO 0);
		F:		OUT	STD_LOGIC_VECTOR(31 DOWNTO 0);
		H:		OUT	STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE DATAFLOW OF EXCEPTIONS IS

COMPONENT IS_NAN IS
	PORT(
		I:	IN	STD_LOGIC_VECTOR(30 DOWNTO 0);
		O:	OUT	STD_LOGIC
	);
END COMPONENT;

COMPONENT IS_ZERO IS
	PORT(
		I:	IN	STD_LOGIC_VECTOR(30 DOWNTO 0);
		O:	OUT	STD_LOGIC
	);
END COMPONENT;

COMPONENT IS_INFINITY IS
	PORT(
		I:	IN	STD_LOGIC_VECTOR(30 DOWNTO 0);
		O:	OUT	STD_LOGIC
	);
END COMPONENT;

COMPONENT OR_C IS
	PORT(
		X:	IN	STD_LOGIC;
		Y:	IN	STD_LOGIC;
		Z:	OUT	STD_LOGIC
	);
END COMPONENT;

COMPONENT XOR_C IS
	PORT(
		X:		IN		STD_LOGIC;
		Y:		IN		STD_LOGIC;
		Z:		OUT		STD_LOGIC
	);
END COMPONENT;

COMPONENT MUX_2_TO_1_32_BITS IS
	PORT(
		SEL:	IN	STD_LOGIC;
		I_0:	IN	STD_LOGIC_VECTOR(31 DOWNTO 0);
		I_1:	IN	STD_LOGIC_VECTOR(31 DOWNTO 0);
		O:		OUT	STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT OR_C_4_BITS IS
	PORT(
		I:	IN	STD_LOGIC_VECTOR(3 DOWNTO 0);
		O:	OUT	STD_LOGIC
	);
END COMPONENT;

COMPONENT FUNCTION_E IS
	PORT(
		N, I, S, O, SI:	IN	STD_LOGIC;
		R:				IN	STD_LOGIC_VECTOR(1 DOWNTO 0);
		F:				OUT	STD_LOGIC_VECTOR(31 DOWNTO 0);
		H:				OUT	STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

SIGNAL O_0, O_1, O_2, O_3, O_4, O_5: STD_LOGIC;
SIGNAL O_6, O_7, O_8: STD_LOGIC;
SIGNAL O_9, O_10: 	STD_LOGIC;
SIGNAL O_11, O_12: 	STD_LOGIC;
SIGNAL O_13: 		STD_LOGIC;
SIGNAL O_14: 		STD_LOGIC;
SIGNAL O_F:			STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL O_H:			STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL P_F:			STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL OR_S:		STD_LOGIC_VECTOR(3 DOWNTO 0);

BEGIN
	
	NAN1:	IS_NAN PORT MAP(B(30 DOWNTO 0), O_0);
	NAN2:	IS_NAN PORT MAP(A(30 DOWNTO 0), O_1);
	ZERO1:	IS_ZERO PORT MAP(A(30 DOWNTO 0), O_2);
	INFI1:	IS_INFINITY PORT MAP(B(30 DOWNTO 0), O_3);
	ZERO2:	IS_ZERO PORT MAP(B(30 DOWNTO 0), O_4);
	INFI2:	IS_INFINITY PORT MAP(A(30 DOWNTO 0), O_5);
	
	OR1:	OR_C PORT MAP(O_0, O_1, O_6);
	OR2:	OR_C PORT MAP(O_2, O_3, O_7);
	OR3:	OR_C PORT MAP(O_4, O_5, O_8);
	
	OR4:	OR_C PORT MAP(O_7, O_8, O_9);
	OR5:	OR_C PORT MAP(O_2, O_4, O_10);
	
	ZERO3:	IS_ZERO PORT MAP(C(30 DOWNTO 0),  O_11);
	INFI3:	IS_INFINITY PORT MAP(C(30 DOWNTO 0), O_12);
	
	XOR1:	XOR_C PORT MAP(O_11, O_10, O_13);
	
	F1:		FUNCTION_E PORT MAP(O_6, O_9, O_13, O_12, C(31), R, O_F, O_H);
	
	OR6:	OR_C_4_BITS PORT MAP(O_H, O_14);
	
	MUX:	MUX_2_TO_1_32_BITS PORT MAP(O_14, C, O_F, P_F);
	
	F <= P_F;
	H <= O_H;
	
END ARCHITECTURE;
