----------------------------------------------------------
--	AUTOR: ULISES MARTINEZ RODRIGUEZ
--	DATE: 2020-11-29
--	DESCRIPTION: REALIZA EL DESPLAZAMIENTO DE 1 BIT A
--				LA DERECHA
----------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY BITSHIFT_RIGHT_96_BITS IS
	PORT(
		A:	IN	STD_LOGIC_VECTOR(95 DOWNTO 0);
		O:	OUT	STD_LOGIC_VECTOR(95 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE DATAFLOW OF BITSHIFT_RIGHT_96_BITS IS
BEGIN
	O(95) <= '0';
	O(94 DOWNTO 0) <= A(95 DOWNTO 1);
END ARCHITECTURE;