----------------------------------------------------------
--	AUTOR: ULISES MARTINEZ RODRIGUEZ
--	DATE: 2020-11-26
--	DESCRIPTION: SUMADOR DE 24 BITS
----------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ADD_24_BITS IS
	PORT(
		CARRYIN:	IN	STD_LOGIC;
		ADDEND1:	IN	STD_LOGIC_VECTOR(23 DOWNTO 0);
		ADDEND2:	IN	STD_LOGIC_VECTOR(23 DOWNTO 0);
		SUM:		OUT	STD_LOGIC_VECTOR(23 DOWNTO 0);
		CARRYOUT:	OUT	STD_LOGIC
	);
END ENTITY;

ARCHITECTURE STRUCTURE OF ADD_24_BITS IS

COMPONENT ADD_8_BITS IS
	PORT(
		CARRYIN:	IN	STD_LOGIC;
		ADDEND1:	IN	STD_LOGIC_VECTOR(7 DOWNTO 0);
		ADDEND2:	IN	STD_LOGIC_VECTOR(7 DOWNTO 0);
		SUM:		OUT	STD_LOGIC_VECTOR(7 DOWNTO 0);
		CARRYOUT:	OUT	STD_LOGIC
	);
END COMPONENT;

SIGNAL	CARRIES:		STD_LOGIC_VECTOR(1 DOWNTO 0);

BEGIN
	
	BITS7DOWNTO0:	ADD_8_BITS PORT MAP(CARRYIN, 	ADDEND1(7 DOWNTO 0),   ADDEND2(7 DOWNTO 0),   SUM(7 DOWNTO 0),   CARRIES(0));
	BITS15DOWNTO8:	ADD_8_BITS PORT MAP(CARRIES(0), ADDEND1(15 DOWNTO 8),  ADDEND2(15 DOWNTO 8),  SUM(15 DOWNTO 8),  CARRIES(1));
	BITS23DOWNTO16:	ADD_8_BITS PORT MAP(CARRIES(1), ADDEND1(23 DOWNTO 16), ADDEND2(23 DOWNTO 16), SUM(23 DOWNTO 16), CARRYOUT);
	

END ARCHITECTURE;