----------------------------------------------------------
--	AUTOR: ULISES MARTINEZ RODRIGUEZ
--	DATE: 2020-12-07
--	DESCRIPTION: DETERMINA SI ES UN NAN
----------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY IS_NAN IS
	PORT(
		I:	IN	STD_LOGIC_VECTOR(30 DOWNTO 0);
		O:	OUT	STD_LOGIC
	);
END ENTITY;

ARCHITECTURE DATAFLOW OF IS_NAN IS
SIGNAL A:	STD_LOGIC;
BEGIN
	A <= I(22) OR I(21) OR I(20) OR I(19) OR I(18) OR I(17) OR I(16) OR I(15) OR I(14) OR I(13)OR I(12) OR I(11) OR I(10) OR I(9) OR I(8) OR I(7) OR I(6) OR I(5) OR I(4) OR I(3) OR I(2) OR I(1) OR I(0);
	O <= '1' WHEN I(30 DOWNTO 23)="11111111" AND A='1' ELSE '0';
END ARCHITECTURE;