----------------------------------------------------------
--	AUTOR: ULISES MARTINEZ RODRIGUEZ
--	DATE: 2020-11-26
--	DESCRIPTION: MULTIPLICADOR DE 24 BITS
----------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MULT_24_BITS IS
	PORT(
		MULTIPLICAND:	IN	STD_LOGIC_VECTOR(23 DOWNTO 0);
		MULTIPLIER:		IN	STD_LOGIC_VECTOR(23 DOWNTO 0);
		PRODUCTHIGH:	OUT	STD_LOGIC_VECTOR(23 DOWNTO 0);
		PRODUCTLOW:		OUT	STD_LOGIC_VECTOR(23 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE STRUCTURE OF MULT_24_BITS IS

COMPONENT ADD_24_BITS IS
	PORT(
		CARRYIN:	IN	STD_LOGIC;
		ADDEND1:	IN	STD_LOGIC_VECTOR(23 DOWNTO 0);
		ADDEND2:	IN	STD_LOGIC_VECTOR(23 DOWNTO 0);
		SUM:		OUT	STD_LOGIC_VECTOR(23 DOWNTO 0);
		CARRYOUT:	OUT	STD_LOGIC
	);
END COMPONENT;

SIGNAL PREPRODUCTS:		STD_LOGIC_VECTOR(575 DOWNTO 0);
SIGNAL PARTIALSADDS:	STD_LOGIC_VECTOR(574 DOWNTO 0);

BEGIN
	
	PREPRODUCT: PROCESS(MULTIPLICAND, MULTIPLIER)
	BEGIN
		FOR J IN 0 TO 23 LOOP
			IF MULTIPLIER(J) = '1' THEN
				PREPRODUCTS((J*24)+23 DOWNTO (J*24)) <= MULTIPLICAND;
			ELSE
				PREPRODUCTS((J*24)+23 DOWNTO (J*24)) <= (OTHERS=>'0');
			END IF;
		END LOOP;
	END PROCESS;
	
	PRODUCTLOW(0)	<= PREPRODUCTS(0);
	ADD0AND1:		ADD_24_BITS PORT MAP('0', '0' & PREPRODUCTS(23 DOWNTO 1), PREPRODUCTS(47 DOWNTO 24), PARTIALSADDS(23 DOWNTO 0), PARTIALSADDS(24));
	
	PRODUCTLOW(1)	<= PARTIALSADDS(0);
	ADD1AND2:	  	ADD_24_BITS PORT MAP('0', PARTIALSADDS(24 DOWNTO 1), PREPRODUCTS(71 DOWNTO 48), PARTIALSADDS(48 DOWNTO 25), PARTIALSADDS(49));
	PRODUCTLOW(2)	<= PARTIALSADDS(25);
	ADD2AND3:	  	ADD_24_BITS PORT MAP('0', PARTIALSADDS(49 DOWNTO 26), PREPRODUCTS(95 DOWNTO 72), PARTIALSADDS(73 DOWNTO 50), PARTIALSADDS(74));
	PRODUCTLOW(3)	<= PARTIALSADDS(50);
	ADD3AND4:	  	ADD_24_BITS PORT MAP('0', PARTIALSADDS(74 DOWNTO 51), PREPRODUCTS(119 DOWNTO 96), PARTIALSADDS(98 DOWNTO 75), PARTIALSADDS(99));
	PRODUCTLOW(4)	<= PARTIALSADDS(75);
	ADD4AND5:	  	ADD_24_BITS PORT MAP('0', PARTIALSADDS(99 DOWNTO 76), PREPRODUCTS(143 DOWNTO 120), PARTIALSADDS(123 DOWNTO 100), PARTIALSADDS(124));
	PRODUCTLOW(5)	<= PARTIALSADDS(100);
	ADD5AND6:	  	ADD_24_BITS PORT MAP('0', PARTIALSADDS(124 DOWNTO 101), PREPRODUCTS(167 DOWNTO 144), PARTIALSADDS(148 DOWNTO 125), PARTIALSADDS(149));
	PRODUCTLOW(6)	<= PARTIALSADDS(125);
	ADD6AND7:	  	ADD_24_BITS PORT MAP('0', PARTIALSADDS(149 DOWNTO 126), PREPRODUCTS(191 DOWNTO 168), PARTIALSADDS(173 DOWNTO 150), PARTIALSADDS(174));
	PRODUCTLOW(7)	<= PARTIALSADDS(150);
	ADD7AND8:	  	ADD_24_BITS PORT MAP('0', PARTIALSADDS(174 DOWNTO 151), PREPRODUCTS(215 DOWNTO 192), PARTIALSADDS(198 DOWNTO 175), PARTIALSADDS(199));
	PRODUCTLOW(8)	<= PARTIALSADDS(175);
	ADD8AND9:	  	ADD_24_BITS PORT MAP('0', PARTIALSADDS(199 DOWNTO 176), PREPRODUCTS(239 DOWNTO 216), PARTIALSADDS(223 DOWNTO 200), PARTIALSADDS(224));
	PRODUCTLOW(9)	<= PARTIALSADDS(200);
	ADD9AND10:	  	ADD_24_BITS PORT MAP('0', PARTIALSADDS(224 DOWNTO 201), PREPRODUCTS(263 DOWNTO 240), PARTIALSADDS(248 DOWNTO 225), PARTIALSADDS(249));
	PRODUCTLOW(10)	<= PARTIALSADDS(225);
	ADD10AND11:	  	ADD_24_BITS PORT MAP('0', PARTIALSADDS(249 DOWNTO 226), PREPRODUCTS(287 DOWNTO 264), PARTIALSADDS(273 DOWNTO 250), PARTIALSADDS(274));
	PRODUCTLOW(11)	<= PARTIALSADDS(250);
	ADD11AND12:	  	ADD_24_BITS PORT MAP('0', PARTIALSADDS(274 DOWNTO 251), PREPRODUCTS(311 DOWNTO 288), PARTIALSADDS(298 DOWNTO 275), PARTIALSADDS(299));
	PRODUCTLOW(12)	<= PARTIALSADDS(275);
	ADD12AND13:	  	ADD_24_BITS PORT MAP('0', PARTIALSADDS(299 DOWNTO 276), PREPRODUCTS(335 DOWNTO 312), PARTIALSADDS(323 DOWNTO 300), PARTIALSADDS(324));
	PRODUCTLOW(13)	<= PARTIALSADDS(300);
	ADD13AND14:	  	ADD_24_BITS PORT MAP('0', PARTIALSADDS(324 DOWNTO 301), PREPRODUCTS(359 DOWNTO 336), PARTIALSADDS(348 DOWNTO 325), PARTIALSADDS(349));
	PRODUCTLOW(14)	<= PARTIALSADDS(325);
	ADD14AND15:	  	ADD_24_BITS PORT MAP('0', PARTIALSADDS(349 DOWNTO 326), PREPRODUCTS(383 DOWNTO 360), PARTIALSADDS(373 DOWNTO 350), PARTIALSADDS(374));
	PRODUCTLOW(15)	<= PARTIALSADDS(350);
	ADD15AND16:	  	ADD_24_BITS PORT MAP('0', PARTIALSADDS(374 DOWNTO 351), PREPRODUCTS(407 DOWNTO 384), PARTIALSADDS(398 DOWNTO 375), PARTIALSADDS(399));
	PRODUCTLOW(16)	<= PARTIALSADDS(375);
	ADD16AND17:	  	ADD_24_BITS PORT MAP('0', PARTIALSADDS(399 DOWNTO 376), PREPRODUCTS(431 DOWNTO 408), PARTIALSADDS(423 DOWNTO 400), PARTIALSADDS(424));
	PRODUCTLOW(17)	<= PARTIALSADDS(400);
	ADD17AND18:	  	ADD_24_BITS PORT MAP('0', PARTIALSADDS(424 DOWNTO 401), PREPRODUCTS(455 DOWNTO 432), PARTIALSADDS(448 DOWNTO 425), PARTIALSADDS(449));
	PRODUCTLOW(18)	<= PARTIALSADDS(425);
	ADD18AND19:	  	ADD_24_BITS PORT MAP('0', PARTIALSADDS(449 DOWNTO 426), PREPRODUCTS(479 DOWNTO 456), PARTIALSADDS(473 DOWNTO 450), PARTIALSADDS(474));
	PRODUCTLOW(19)	<= PARTIALSADDS(450);
	ADD19AND20:	  	ADD_24_BITS PORT MAP('0', PARTIALSADDS(474 DOWNTO 451), PREPRODUCTS(503 DOWNTO 480), PARTIALSADDS(498 DOWNTO 475), PARTIALSADDS(499));
	PRODUCTLOW(20)	<= PARTIALSADDS(475);
	ADD20AND21:	  	ADD_24_BITS PORT MAP('0', PARTIALSADDS(499 DOWNTO 476), PREPRODUCTS(527 DOWNTO 504), PARTIALSADDS(523 DOWNTO 500), PARTIALSADDS(524));
	PRODUCTLOW(21)	<= PARTIALSADDS(500);
	ADD21AND22:	  	ADD_24_BITS PORT MAP('0', PARTIALSADDS(524 DOWNTO 501), PREPRODUCTS(551 DOWNTO 528), PARTIALSADDS(548 DOWNTO 525), PARTIALSADDS(549));
	PRODUCTLOW(22)	<= PARTIALSADDS(525);
	ADD22AND23:	  	ADD_24_BITS PORT MAP('0', PARTIALSADDS(549 DOWNTO 526), PREPRODUCTS(575 DOWNTO 552), PARTIALSADDS(573 DOWNTO 550), PARTIALSADDS(574));	
	
	PRODUCTLOW(23)	<= PARTIALSADDS(550);
	PRODUCTHIGH		<= PARTIALSADDS(574 DOWNTO 551);
	
END ARCHITECTURE;